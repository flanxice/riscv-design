`timescale 1ns / 1ps
module Risc5CPU(
    input clk,
    input reset,
    output[1:0] JumpFlag,
    output [31:0] Instruction_id,
    output [31:0] ALU_A,
    output [31:0] ALU_B,
    output [31:0] ALUResult_ex,
    output [31:0] PC,
    output [31:0] MemDout_mem,
    output Stall);

wire IFWrite, IF_flush;
wire [31:0] JumpAddr;
wire [31:0] Instruction_if, PC;
IF IF_STATE(.clk(clk), .reset(reset), .Branch(JumpFlag[0]), .Jump(JumpFlag[1]),
    .IFWrite(IFWrite), .JumpAddr(JumpAddr), .Instruction_if(Instruction_if),
    .PC(PC), .IF_flush(IF_flush));

wire [31:0] Instruction_id, PC_id;
IF_ID_PipeReg PR1(.clk(clk), .EN(IFWrite), .R((IF_flush | reset)),
    .PC_in_c(PC), .Instruction_in_c(Instruction_if),
    .PC_out_c(PC_id), .Instruction_out_c(Instruction_id));

wire RegWrite_wb, MemtoReg_id, RegWrite_id, MemWrite_id, MemRead_id, ALUSrcA_id;   
wire [4:0] rdAddr_ex, rs1Addr_id, rs2Addr_id, rdAddr_id;
wire [31:0] RegWriteData_wb, Imm_id, rs1Data_id, rs2Data_id;
wire [3:0] ALUCode_id;
wire [1:0] ALUSrcB_id;
ID ID_STATE(.clk(clk), .Instruction_id(Instruction_id), .PC_id(PC_id),
    .RegWrite_wb(RegWrite_wb), .rdAddr_wb(rdAddr_wb), .RegWriteData_wb(RegWriteData_wb),
    .MemRead_ex(MemRead_ex), .rdAddr_ex(rdAddr_ex), .MemtoReg_id(MemtoReg_id),
    .RegWrite_id(RegWrite_id), .MemWrite_id(MemWrite_id),
    .MemRead_id(MemRead_id), .ALUCode_id(ALUCode_id), .ALUSrcA_id(ALUSrcA_id),
    .ALUSrcB_id(ALUSrcB_id), .Stall(Stall), .Branch(JumpFlag[0]), .Jump(JumpFlag[1]),
    .IFWrite(IFWrite), .JumpAddr(JumpAddr), .Imm_id(Imm_id),
    .rs1Data_id(rs1Data_id), .rs2Data_id(rs2Data_id),
	.rs1Addr_id(rs1Addr_id), .rs2Addr_id(rs2Addr_id), .rdAddr_id(rdAddr_id));

wire MemtoReg_ex, RegWrite_ex, MemWrite_ex, MemRead_ex, ALUSrcA_ex;
wire [3:0] ALUCode_ex;
wire [1:0] ALUSrcB_ex;
wire [4:0] rs1Addr_ex, rs2Addr_ex;
wire [31:0] PC_ex, rs1Data_ex, rs2Data_ex, Imm_ex;
ID_EX_PipeReg PR2(.clk(clk), .R(Stall | reset), .MemtoReg_id(MemtoReg_id), .RegWrite_id(RegWrite_id), 
    .MemWrite_id(MemWrite_id), .MemRead_id(MemRead_id), .ALUCode_id(ALUCode_id),
    .ALUSrcA_id(ALUSrcA_id), .ALUSrcB_id(ALUSrcB_id), .rs1Addr_id(rs1Addr_id), .rs2Addr_id(rs2Addr_id), .rdAddr_id(rdAddr_id),
    .PC_id(PC_id), .rs1Data_id(rs1Data_id), .rs2Data_id(rs2Data_id),
    .Imm_id(Imm_id), .MemtoReg_ex(MemtoReg_ex), .RegWrite_ex(RegWrite_ex), .MemWrite_ex(MemWrite_ex), .MemRead_ex(MemRead_ex),
    .ALUCode_ex(ALUCode_ex), .ALUSrcA_ex(ALUSrcA_ex), .ALUSrcB_ex(ALUSrcB_ex),
    .rdAddr_ex(rdAddr_ex), .rs1Addr_ex(rs1Addr_ex), .rs2Addr_ex(rs2Addr_ex),
    .PC_ex(PC_ex), .rs1Data_ex(rs1Data_ex), .rs2Data_ex(rs2Data_ex), .Imm_ex(Imm_ex));

wire [31:0] ALUResult_mem, ALUResult_ex, MemWriteData_ex;
wire [4:0] rdAddr_mem, rdAddr_wb;
wire RegWrite_mem, RegWrite_wb;
EX EX_STATE(.ALUCode_ex(ALUCode_ex), .ALUSrcA_ex(ALUSrcA_ex), .ALUSrcB_ex(ALUSrcB_ex),
    .Imm_ex(Imm_ex), .rs1Addr_ex(rs1Addr_ex), .rs2Addr_ex(rs2Addr_ex), .rs1Data_ex(rs1Data_ex),
    .rs2Data_ex(rs2Data_ex), .PC_ex(PC_ex), .RegWriteData_wb(RegWriteData_wb),
    .ALUResult_mem(ALUResult_mem), .rdAddr_mem(rdAddr_mem), .rdAddr_wb(rdAddr_wb),
    .RegWrite_mem(RegWrite_mem), .RegWrite_wb(RegWrite_wb), .ALUResult_ex(ALUResult_ex),
    .MemWriteData_ex(MemWriteData_ex), .ALU_A(ALU_A), .ALU_B(ALU_B));

wire MemtoReg_mem, RegWrite_mem, MemWrite_mem;
wire [31:0] MemWriteData_mem;
EX_mem_PinpeReg PR3(.clk(clk), .MemtoReg_ex(MemtoReg_ex), .RegWrite_ex(RegWrite_ex), .MemWrite_ex(MemWrite_ex),
    .ALUout(ALUResult_ex), .MemWriteData_ex(MemWriteData_ex), .rdAddr_ex(rdAddr_ex), 
    .MemtoReg_mem(MemtoReg_mem), .RegWrite_mem(RegWrite_mem), .MemWrite_mem(MemWrite_mem),
    .ALUResult_mem(ALUResult_mem), .MemWriteData_mem(MemWriteData_mem), .rdAddr_mem(rdAddr_mem));

DRAM DRAM0(.a(ALUResult_mem[7:2]), .d(MemWriteData_mem), .clk(clk),
    .we(MemWrite_mem), .spo(MemDout_mem));

wire MemtoReg_wb, RegWrite_wb;
wire [31:0] MemDout_wb, ALUResult_wb;
DM_WB_PipeReg PR4(
.clk(clk), .MemtoReg_mem(MemtoReg_mem), .RegWrite_mem(RegWrite_mem),
.MemDout_mem(MemDout_mem), .ALUResult_mem(ALUResult_mem),
.rdAddr_mem(rdAddr_mem), .MemtoReg_wb(MemtoReg_wb), .RegWrite_wb(RegWrite_wb),
.MemDout_wb(MemDout_wb), .ALUResult_wb(ALUResult_wb), .rdAddr_wb(rdAddr_wb));

WB WB_STATE(
    .MemtoReg_wb(MemtoReg_wb), .MemDout_wb(MemDout_wb), .ALUResult_wb(ALUResult_wb),
    .RegWriteData_wb(RegWriteData_wb));

endmodule
